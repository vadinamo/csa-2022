`ifndef SWORD
`define SWORD

package sword;
	typedef enum logic [1:0] {S0, S1} sword_state;
endpackage

`endif