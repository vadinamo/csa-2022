module fulladder(input logic a, b, cin,
										output logic sum)