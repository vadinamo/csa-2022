module testbench(); 
	logic clk, reset;
	logic n, s, w, e, win, lose;
	logic [1:0] expected;
	logic [31:0] vectornum, errors;
	logic [7:0] testvectors[10000:0];
	logic r;
	
	task2 dut(clk, reset, n, s, w, e, win, lose);
	
	always
		begin
			clk=1; #5; clk=0; #5; 
		end
		
	initial
		begin
			$readmemb("test.tv", testvectors); 
			vectornum = 0; errors = 0; reset = 1; #22; reset = 0; 
		end
		
	always @(posedge clk) 
		begin
			#1; {r, n, s, w, e, expected} = testvectors[vectornum];
			if(r)
				begin
					reset = 1; #22; reset = 0;
				end
		end
		
	always @(negedge clk) 
		if (~reset) begin
			if ({win, lose} !== expected) begin
				$display("Error: inputs = %b", {reset, n, s, w, e});
				$display(" outputs = %b %b (%b expected)", win, lose, expected); 
				errors = errors + 1; 
			end
			vectornum = vectornum + 1;
			if (testvectors[vectornum] === 8'bx) begin
				$display("%d tests completed with %d errors", vectornum, errors); 
				$stop; 
			end
		end
endmodule