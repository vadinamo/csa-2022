`ifndef TREASURE
`define TREASURE

package treasure;
	typedef enum logic [1:0] {T0, T1} treasure_state;
endpackage

`endif