`ifndef ROOMS
`define ROOMS

package rooms;
	typedef enum logic [3:0] {R1, R2, R3, R4, R5, R6, R7, R8, R9} room_states;
endpackage

`endif